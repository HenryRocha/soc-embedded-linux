
module niosLab2 (
	clk_clk,
	reset_reset_n,
	leds_leds,
	buts_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	leds_leds;
	input	[3:0]	buts_export;
endmodule
